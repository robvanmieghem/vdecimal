module vdecimal

fn test_ci() ? {
}
